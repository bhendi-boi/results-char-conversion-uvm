class rcc_configuration extends uvm_object;
  `uvm_object_utils(rcc_configuration)

  function new(string name = "");
    super.new(name);
  endfunction : new

endclass : rcc_configuration
